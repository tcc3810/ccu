`include "FA.v"
`include "HA.v"
module MPY(clk, a, b, p);
    input clk;
    input [31:0] a, b;
    output [63:0] p;
    wire [32:0] add0, add1, add2, add3, add4, add5, add6, add7, add8, add9, 
				add10, add11, add12, add13, add14, add15, add16, add17, add18, add19, 
				add20, add21, add22, add23, add24, add25, add26, add27, add28, add29, add30, add31;
    wire [63:0] add0_ext;
    wire [62:0] add1_ext;
    wire [61:0] add2_ext;
	wire [60:0] add3_ext;
	wire [59:0] add4_ext;
	wire [58:0] add5_ext;
	wire [57:0] add6_ext;
	wire [56:0] add7_ext;
	wire [55:0] add8_ext;
	wire [54:0] add9_ext;
	wire [53:0] add10_ext;
	wire [52:0] add11_ext;
	wire [51:0] add12_ext;
	wire [50:0] add13_ext;
	wire [49:0] add14_ext;
	wire [48:0] add15_ext;
	wire [47:0] add16_ext;
	wire [46:0] add17_ext;
	wire [45:0] add18_ext;
	wire [44:0] add19_ext;
	wire [43:0] add20_ext;
	wire [42:0] add21_ext;
	wire [41:0] add22_ext;
	wire [40:0] add23_ext;
	wire [39:0] add24_ext;
	wire [38:0] add25_ext;
	wire [37:0] add26_ext;
	wire [36:0] add27_ext;
	wire [35:0] add28_ext;
	wire [34:0] add29_ext;
	wire [33:0] add30_ext;
	
    wire [62:0] s0;
    wire [61:0] s1;
    wire [60:0] s2;
	wire [59:0] s3;
	wire [58:0] s4;
	wire [57:0] s5;
	wire [56:0] s6;
	wire [55:0] s7;
	wire [54:0] s8;
	wire [53:0] s9;
	wire [52:0] s10;
	wire [51:0] s11;
	wire [50:0] s12;
	wire [49:0] s13;
	wire [48:0] s14;
	wire [47:0] s15;
	wire [46:0] s16;
	wire [45:0] s17;
	wire [44:0] s18;
	wire [43:0] s19;
	wire [42:0] s20;
	wire [41:0] s21;
	wire [40:0] s22;
	wire [39:0] s23;
	wire [38:0] s24;
	wire [37:0] s25;
	wire [36:0] s26;
	wire [35:0] s27;
	wire [34:0] s28;
	wire [33:0] s29;
	wire [32:0] s30;
	
    booth_add booth1(a, {b[0],1'b0}, add0);
    booth_add booth2(a, b[1:0], add1);
    booth_add booth3(a, b[2:1], add2);
    booth_add booth4(a, b[3:2], add3);
	booth_add booth5(a, b[4:3], add4);
	booth_add booth6(a, b[5:4], add5);
	booth_add booth7(a, b[6:5], add6);
	booth_add booth8(a, b[7:6], add7);
	booth_add booth9(a, b[8:7], add8);
	booth_add booth10(a, b[9:8], add9);
	booth_add booth11(a, b[10:9], add10);
	booth_add booth12(a, b[11:10], add11);
	booth_add booth13(a, b[12:11], add12);
	booth_add booth14(a, b[13:12], add13);
	booth_add booth15(a, b[14:13], add14);
	booth_add booth16(a, b[15:14], add15);
	booth_add booth17(a, b[16:15], add16);
	booth_add booth18(a, b[17:16], add17);
	booth_add booth19(a, b[18:17], add18);
	booth_add booth20(a, b[19:18], add19);
	booth_add booth21(a, b[20:19], add20);
	booth_add booth22(a, b[21:20], add21);
	booth_add booth23(a, b[22:21], add22);
	booth_add booth24(a, b[23:22], add23);
	booth_add booth25(a, b[24:23], add24);
	booth_add booth26(a, b[25:24], add25);
	booth_add booth27(a, b[26:25], add26);
	booth_add booth28(a, b[27:26], add27);
	booth_add booth29(a, b[28:27], add28);
	booth_add booth30(a, b[29:28], add29);
	booth_add booth31(a, b[30:29], add30);
	booth_add booth32(a, b[31:30], add31);
	
    assign add0_ext = {{31{add0[32]}},add0};
    assign add1_ext = {{30{add1[32]}},add1};
    assign add2_ext = {{29{add2[32]}},add2};
	assign add3_ext = {{28{add3[32]}},add3};
    assign add4_ext = {{27{add4[32]}},add4};
    assign add5_ext = {{26{add5[32]}},add5};
	assign add6_ext = {{25{add6[32]}},add6};
    assign add7_ext = {{24{add7[32]}},add7};
    assign add8_ext = {{23{add8[32]}},add8};
	assign add9_ext = {{22{add9[32]}},add9};
    assign add10_ext = {{21{add10[32]}},add10};
    assign add11_ext = {{20{add11[32]}},add11};
	assign add12_ext = {{19{add12[32]}},add12};
    assign add13_ext = {{18{add13[32]}},add13};
    assign add14_ext = {{17{add14[32]}},add14};
	assign add15_ext = {{16{add15[32]}},add15};
    assign add16_ext = {{15{add16[32]}},add16};
    assign add17_ext = {{14{add17[32]}},add17};
	assign add18_ext = {{13{add18[32]}},add18};
    assign add19_ext = {{12{add19[32]}},add19};
    assign add20_ext = {{11{add20[32]}},add20};
	assign add21_ext = {{10{add21[32]}},add21};
    assign add22_ext = {{9{add22[32]}},add22};
    assign add23_ext = {{8{add23[32]}},add23};
	assign add24_ext = {{7{add24[32]}},add24};
    assign add25_ext = {{6{add25[32]}},add25};
    assign add26_ext = {{5{add26[32]}},add26};
	assign add27_ext = {{4{add27[32]}},add27};
	assign add28_ext = {{3{add28[32]}},add28};
	assign add29_ext = {{2{add29[32]}},add29};
	assign add30_ext = {add30[32],add30};
	
    HA1FA62 HA1FA62_u1(clk, add0_ext[63:1], add1_ext, s0);
    HA1FA61 HA1FA61_u1(clk, s0[62:1], add2_ext, s1);
    HA1FA60 HA1FA60_u1(clk, s1[61:1], add3_ext, s2);
	HA1FA59 HA1FA59_u1(clk, s2[60:1], add4_ext, s3);
	HA1FA58 HA1FA58_u1(clk, s3[59:1], add5_ext, s4);
	HA1FA57 HA1FA57_u1(clk, s4[58:1], add6_ext, s5);
	HA1FA56 HA1FA56_u1(clk, s5[57:1], add7_ext, s6);
	HA1FA55 HA1FA55_u1(clk, s6[56:1], add8_ext, s7);
	HA1FA54 HA1FA54_u1(clk, s7[55:1], add9_ext, s8);
	HA1FA53 HA1FA53_u1(clk, s8[54:1], add10_ext, s9);
	HA1FA52 HA1FA52_u1(clk, s9[53:1], add11_ext, s10);
	HA1FA51 HA1FA51_u1(clk, s10[52:1], add12_ext, s11);
	HA1FA50 HA1FA50_u1(clk, s11[51:1], add13_ext, s12);
	HA1FA49 HA1FA49_u1(clk, s12[50:1], add14_ext, s13);
	HA1FA48 HA1FA48_u1(clk, s13[49:1], add15_ext, s14);
	HA1FA47 HA1FA47_u1(clk, s14[48:1], add16_ext, s15);
	HA1FA46 HA1FA46_u1(clk, s15[47:1], add17_ext, s16);
	HA1FA45 HA1FA45_u1(clk, s16[46:1], add18_ext, s17);
	HA1FA44 HA1FA44_u1(clk, s17[45:1], add19_ext, s18);
	HA1FA43 HA1FA43_u1(clk, s18[44:1], add20_ext, s19);
	HA1FA42 HA1FA42_u1(clk, s19[43:1], add21_ext, s20);
	HA1FA41 HA1FA41_u1(clk, s20[42:1], add22_ext, s21);
	HA1FA40 HA1FA40_u1(clk, s21[41:1], add23_ext, s22);
	HA1FA39 HA1FA39_u1(clk, s22[40:1], add24_ext, s23);
	HA1FA38 HA1FA38_u1(clk, s23[39:1], add25_ext, s24);
	HA1FA37 HA1FA37_u1(clk, s24[38:1], add26_ext, s25);
	HA1FA36 HA1FA36_u1(clk, s25[37:1], add27_ext, s26);
	HA1FA35 HA1FA35_u1(clk, s26[36:1], add28_ext, s27);
	HA1FA34 HA1FA34_u1(clk, s27[35:1], add29_ext, s28);
	HA1FA33 HA1FA33_u1(clk, s28[34:1], add30_ext, s29);
	HA1FA32 HA1FA32_u1(clk, s29[33:1], add31, s30);
	
    assign p[0] = add0_ext[0];
    assign p[1] = s0[0];
    assign p[2] = s1[0];
	assign p[3] = s2[0];
	assign p[4] = s3[0];
	assign p[5] = s4[0];
	assign p[6] = s5[0];
	assign p[7] = s6[0];
	assign p[8] = s7[0];
	assign p[9] = s8[0];
	assign p[10] = s9[0];
	assign p[11] = s10[0];
	assign p[12] = s11[0];
	assign p[13] = s12[0];
	assign p[14] = s13[0];
	assign p[15] = s14[0];
	assign p[16] = s15[0];
	assign p[17] = s16[0];
	assign p[18] = s17[0];
	assign p[19] = s18[0];
	assign p[20] = s19[0];
	assign p[21] = s20[0];
	assign p[22] = s21[0];
	assign p[23] = s22[0];
	assign p[24] = s23[0];
	assign p[25] = s24[0];
	assign p[26] = s25[0];
	assign p[27] = s26[0];
	assign p[28] = s27[0];
	assign p[29] = s28[0];
	assign p[30] = s29[0];
    assign p[63:31] = s30;
endmodule

module booth_add(a, b, ab);
    input [31:0] a;
    input [1:0] b;
    wire signed [32:0] a_ext;
    output [32:0] ab;

    assign a_ext = {a[31],a};
    assign ab = (b==2'b01) ? a_ext:
                (b==2'b10) ? -a_ext:
                             33'b0;                                
endmodule

////////////////////////////////////////////////////////////////////////////////////

module HA1FA32(clk, a, b, s);
    input clk;
    input [32:0] a;
    input [32:0] b;
    output [32:0] s;
	
    wire [32:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);

    assign cout = carry[32];
endmodule

module HA1FA33(clk, a, b, s);
    input clk;
    input [33:0] a;
    input [33:0] b;
    output [33:0] s;
	
    wire [33:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);

    assign cout = carry[33];
endmodule

module HA1FA34(clk, a, b, s);
    input clk;
    input [34:0] a;
    input [34:0] b;
    output [34:0] s;
	
    wire [34:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);

    assign cout = carry[34];
endmodule

module HA1FA35(clk, a, b, s);
    input clk;
    input [35:0] a;
    input [35:0] b;
    output [35:0] s;
	
    wire [35:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);

    assign cout = carry[35];
endmodule

module HA1FA36(clk, a, b, s);
    input clk;
    input [36:0] a;
    input [36:0] b;
    output [36:0] s;
	
    wire [36:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);

    assign cout = carry[36];
endmodule

module HA1FA37(clk, a, b, s);
    input clk;
    input [37:0] a;
    input [37:0] b;
    output [37:0] s;
	
    wire [37:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);

    assign cout = carry[37];
endmodule

module HA1FA38(clk, a, b, s);
    input clk;
    input [38:0] a;
    input [38:0] b;
    output [38:0] s;
	
    wire [38:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);

    assign cout = carry[38];
endmodule

module HA1FA39(clk, a, b, s);
    input clk;
    input [39:0] a;
    input [39:0] b;
    output [39:0] s;
	
    wire [39:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);

    assign cout = carry[39];
endmodule

module HA1FA40(clk, a, b, s);
    input clk;
    input [40:0] a;
    input [40:0] b;
    output [40:0] s;
	
    wire [40:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);

    assign cout = carry[40];
endmodule

module HA1FA41(clk, a, b, s);
    input clk;
    input [41:0] a;
    input [41:0] b;
    output [41:0] s;
	
    wire [41:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);

    assign cout = carry[41];
endmodule

module HA1FA42(clk, a, b, s);
    input clk;
    input [42:0] a;
    input [42:0] b;
    output [42:0] s;
	
    wire [42:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);

    assign cout = carry[42];
endmodule

module HA1FA43(clk, a, b, s);
    input clk;
    input [43:0] a;
    input [43:0] b;
    output [43:0] s;
	
    wire [43:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);

    assign cout = carry[43];
endmodule

module HA1FA44(clk, a, b, s);
    input clk;
    input [44:0] a;
    input [44:0] b;
    output [44:0] s;
	
    wire [44:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);

    assign cout = carry[44];
endmodule

module HA1FA45(clk, a, b, s);
    input clk;
    input [45:0] a;
    input [45:0] b;
    output [45:0] s;
	
    wire [45:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);

    assign cout = carry[45];
endmodule

module HA1FA46(clk, a, b, s);
    input clk;
    input [46:0] a;
    input [46:0] b;
    output [46:0] s;
	
    wire [46:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);

    assign cout = carry[46];
endmodule

module HA1FA47(clk, a, b, s);
    input clk;
    input [47:0] a;
    input [47:0] b;
    output [47:0] s;
	
    wire [47:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);

    assign cout = carry[47];
endmodule

module HA1FA48(clk, a, b, s);
    input clk;
    input [48:0] a;
    input [48:0] b;
    output [48:0] s;
	
    wire [48:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);

    assign cout = carry[48];
endmodule

module HA1FA49(clk, a, b, s);
    input clk;
    input [49:0] a;
    input [49:0] b;
    output [49:0] s;
	
    wire [49:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);

    assign cout = carry[49];
endmodule

module HA1FA50(clk, a, b, s);
    input clk;
    input [50:0] a;
    input [50:0] b;
    output [50:0] s;
	
    wire [50:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);

    assign cout = carry[50];
endmodule

module HA1FA51(clk, a, b, s);
    input clk;
    input [51:0] a;
    input [51:0] b;
    output [51:0] s;
	
    wire [51:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);

    assign cout = carry[51];
endmodule

module HA1FA52(clk, a, b, s);
    input clk;
    input [52:0] a;
    input [52:0] b;
    output [52:0] s;
	
    wire [52:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);

    assign cout = carry[52];
endmodule

module HA1FA53(clk, a, b, s);
    input clk;
    input [53:0] a;
    input [53:0] b;
    output [53:0] s;
	
    wire [53:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);

    assign cout = carry[53];
endmodule

module HA1FA54(clk, a, b, s);
    input clk;
    input [54:0] a;
    input [54:0] b;
    output [54:0] s;
	
    wire [54:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);

    assign cout = carry[54];
endmodule

module HA1FA55(clk, a, b, s);
    input clk;
    input [55:0] a;
    input [55:0] b;
    output [55:0] s;
	
    wire [55:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);

    assign cout = carry[55];
endmodule

module HA1FA56(clk, a, b, s);
    input clk;
    input [56:0] a;
    input [56:0] b;
    output [56:0] s;
	
    wire [56:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);

    assign cout = carry[56];
endmodule

module HA1FA57(clk, a, b, s);
    input clk;
    input [57:0] a;
    input [57:0] b;
    output [57:0] s;
	
    wire [57:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);

    assign cout = carry[57];
endmodule

module HA1FA58(clk, a, b, s);
    input clk;
    input [58:0] a;
    input [58:0] b;
    output [58:0] s;
	
    wire [58:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);
    FA FA58(clk,a[58],b[58],carry[57],s[58],carry[58]);

    assign cout = carry[58];
endmodule

module HA1FA59(clk, a, b, s);
    input clk;
    input [59:0] a;
    input [59:0] b;
    output [59:0] s;
	
    wire [59:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);
    FA FA58(clk,a[58],b[58],carry[57],s[58],carry[58]);
    FA FA59(clk,a[59],b[59],carry[58],s[59],carry[59]);

    assign cout = carry[59];
endmodule

module HA1FA60(clk, a, b, s);
    input clk;
    input [60:0] a;
    input [60:0] b;
    output [60:0] s;
	
    wire [60:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);
    FA FA58(clk,a[58],b[58],carry[57],s[58],carry[58]);
    FA FA59(clk,a[59],b[59],carry[58],s[59],carry[59]);
    FA FA60(clk,a[60],b[60],carry[59],s[60],carry[60]);

    assign cout = carry[60];
endmodule

module HA1FA61(clk, a, b, s);
    input clk;
    input [61:0] a;
    input [61:0] b;
    output [61:0] s;
	
    wire [61:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);
    FA FA58(clk,a[58],b[58],carry[57],s[58],carry[58]);
    FA FA59(clk,a[59],b[59],carry[58],s[59],carry[59]);
    FA FA60(clk,a[60],b[60],carry[59],s[60],carry[60]);
    FA FA61(clk,a[61],b[61],carry[60],s[61],carry[61]);

    assign cout = carry[61];
endmodule

module HA1FA62(clk, a, b, s);
    input clk;
    input [62:0] a;
    input [62:0] b;
    output [62:0] s;
	
    wire [62:0] carry;
    wire cout;
    HA HA1(clk,a[0],b[0],s[0],carry[0]);
    FA FA1(clk,a[1],b[1],carry[0],s[1],carry[1]);
    FA FA2(clk,a[2],b[2],carry[1],s[2],carry[2]);
    FA FA3(clk,a[3],b[3],carry[2],s[3],carry[3]);
    FA FA4(clk,a[4],b[4],carry[3],s[4],carry[4]);
    FA FA5(clk,a[5],b[5],carry[4],s[5],carry[5]);
    FA FA6(clk,a[6],b[6],carry[5],s[6],carry[6]);
    FA FA7(clk,a[7],b[7],carry[6],s[7],carry[7]);
    FA FA8(clk,a[8],b[8],carry[7],s[8],carry[8]);
    FA FA9(clk,a[9],b[9],carry[8],s[9],carry[9]);
    FA FA10(clk,a[10],b[10],carry[9],s[10],carry[10]);
    FA FA11(clk,a[11],b[11],carry[10],s[11],carry[11]);
    FA FA12(clk,a[12],b[12],carry[11],s[12],carry[12]);
    FA FA13(clk,a[13],b[13],carry[12],s[13],carry[13]);
    FA FA14(clk,a[14],b[14],carry[13],s[14],carry[14]);
    FA FA15(clk,a[15],b[15],carry[14],s[15],carry[15]);
    FA FA16(clk,a[16],b[16],carry[15],s[16],carry[16]);
    FA FA17(clk,a[17],b[17],carry[16],s[17],carry[17]);
    FA FA18(clk,a[18],b[18],carry[17],s[18],carry[18]);
    FA FA19(clk,a[19],b[19],carry[18],s[19],carry[19]);
    FA FA20(clk,a[20],b[20],carry[19],s[20],carry[20]);
    FA FA21(clk,a[21],b[21],carry[20],s[21],carry[21]);
    FA FA22(clk,a[22],b[22],carry[21],s[22],carry[22]);
    FA FA23(clk,a[23],b[23],carry[22],s[23],carry[23]);
    FA FA24(clk,a[24],b[24],carry[23],s[24],carry[24]);
    FA FA25(clk,a[25],b[25],carry[24],s[25],carry[25]);
    FA FA26(clk,a[26],b[26],carry[25],s[26],carry[26]);
    FA FA27(clk,a[27],b[27],carry[26],s[27],carry[27]);
    FA FA28(clk,a[28],b[28],carry[27],s[28],carry[28]);
    FA FA29(clk,a[29],b[29],carry[28],s[29],carry[29]);
    FA FA30(clk,a[30],b[30],carry[29],s[30],carry[30]);
    FA FA31(clk,a[31],b[31],carry[30],s[31],carry[31]);
    FA FA32(clk,a[32],b[32],carry[31],s[32],carry[32]);
    FA FA33(clk,a[33],b[33],carry[32],s[33],carry[33]);
    FA FA34(clk,a[34],b[34],carry[33],s[34],carry[34]);
    FA FA35(clk,a[35],b[35],carry[34],s[35],carry[35]);
    FA FA36(clk,a[36],b[36],carry[35],s[36],carry[36]);
    FA FA37(clk,a[37],b[37],carry[36],s[37],carry[37]);
    FA FA38(clk,a[38],b[38],carry[37],s[38],carry[38]);
    FA FA39(clk,a[39],b[39],carry[38],s[39],carry[39]);
    FA FA40(clk,a[40],b[40],carry[39],s[40],carry[40]);
    FA FA41(clk,a[41],b[41],carry[40],s[41],carry[41]);
    FA FA42(clk,a[42],b[42],carry[41],s[42],carry[42]);
    FA FA43(clk,a[43],b[43],carry[42],s[43],carry[43]);
    FA FA44(clk,a[44],b[44],carry[43],s[44],carry[44]);
    FA FA45(clk,a[45],b[45],carry[44],s[45],carry[45]);
    FA FA46(clk,a[46],b[46],carry[45],s[46],carry[46]);
    FA FA47(clk,a[47],b[47],carry[46],s[47],carry[47]);
    FA FA48(clk,a[48],b[48],carry[47],s[48],carry[48]);
    FA FA49(clk,a[49],b[49],carry[48],s[49],carry[49]);
    FA FA50(clk,a[50],b[50],carry[49],s[50],carry[50]);
    FA FA51(clk,a[51],b[51],carry[50],s[51],carry[51]);
    FA FA52(clk,a[52],b[52],carry[51],s[52],carry[52]);
    FA FA53(clk,a[53],b[53],carry[52],s[53],carry[53]);
    FA FA54(clk,a[54],b[54],carry[53],s[54],carry[54]);
    FA FA55(clk,a[55],b[55],carry[54],s[55],carry[55]);
    FA FA56(clk,a[56],b[56],carry[55],s[56],carry[56]);
    FA FA57(clk,a[57],b[57],carry[56],s[57],carry[57]);
    FA FA58(clk,a[58],b[58],carry[57],s[58],carry[58]);
    FA FA59(clk,a[59],b[59],carry[58],s[59],carry[59]);
    FA FA60(clk,a[60],b[60],carry[59],s[60],carry[60]);
    FA FA61(clk,a[61],b[61],carry[60],s[61],carry[61]);
    FA FA62(clk,a[62],b[62],carry[61],s[62],carry[62]);

    assign cout = carry[62];
endmodule
