module lab5_birth(	
		input [2:0] cnt,
		output [3:0] birth_num,
		output reg [6:0] seg_data
	);

//**CODE_CONVERTER**//

/////////////////////


//**BCD_to_7SEG**//

///////////////////
	
endmodule